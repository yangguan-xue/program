module x(
    input wire A,B,C,
    output wire F
);
    assign F = A & C;
endmodule